`default_nettype none

module tt_um_htfab_cells (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

cell_mux cm_inst (
    .page(ui_in[3:0]),
    .in({uio_in[1:0], ui_in[7:4]}),
    .out(uo_out)
);

assign uio_out = 0;
assign uio_oe = 0;
wire _unused = &{ena, clk, rst_n, uio_in[7:2], 1'b0};

endmodule
